`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Copyright: Chris Larsen, 2022
//
// Create Date: 11/07/2022 09:27:02 AM
// Design Name:
// Module Name: recip_x
// Project Name:
// Target Devices:
// Tool Versions:
// Description: Module to compute the reciprocal of a number D.
//              Normally, we want to compute the reciprocal of a divisor so
//              we can avoid floating point division; multiplication by the
//              reciprocal is almost always much faster. And when performing
//              linear algebra the same divisor is often used multiple times
//              for operations such as normalizing a vector.
//
//              In its present form the module is combinatorial logic.
//              Eventually it will need to be a state machine.
//
//              Inputs:
//              - d: The divisor for which we wish to compute the reciprocal.
//              - ra: The rounding attribute to be used when truncating the
//                    result to fit into the final binary16/-32/-64/-128 result.
//              Outputs:
//              - r: The computed reciprocal value.
//              - rFlags: Flags telling the system which type of value (sNaN,
//                qNaN, Infinity, etc.) is being returned by the module.
//              - exception: Exceptions generated by the module.
//
// Dependencies: fp_class.sv
//               ieee-754-flags.vh
//               padder11.v
//               padder24.v
//               PijGij.v
//               round.v
//               X0.v
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module recip_x(d, ra, r, rFlags, exception);
  parameter NEXP = 5;
  parameter NSIG = 10;
  `include "ieee-754-flags.vh"
  localparam CLOG2_NSIG = $clog2(NSIG+1);
  input [NEXP+NSIG:0] d;
  input [NRAS-1:0] ra;
  output [NEXP+NSIG:0] r;
  output [NTYPES-1:0] rFlags;
  reg [NTYPES-1:0] rFlags;
  output [NEXCEPTIONS-1:0] exception;
  reg [NEXCEPTIONS-1:0] exception;

  localparam hNSIG = 10;

  wire inexact, inexactH, inexactX;

  wire signed [NEXP+1:0] dExp, expOut;
  reg signed [NEXP+1:0] rExp, expIn, normExp = 0;
  wire [0:-NSIG] dSigWire, sigOut;
  wire [NTYPES-1:0] dFlags;
  fp_class #(NEXP,NSIG) dClass(d, dExp, dSigWire, dFlags);

  wire [0:-NSIG-1] x0;
  X0 #(NEXP,NSIG) U0(dSigWire[-1:-hNSIG], x0);

  reg [0:-(3*NSIG+2)] sigIn;

  reg [NEXP+NSIG:0] alwaysR;

  reg si;
  integer i;
  always @(*)
    begin
      rFlags = 0;
      exception = 0;

      case (dFlags)
        6'b100000: begin // sNaN
            {alwaysR, rFlags} = {d, dFlags};
          end
        6'b010000: begin // qNaN
            {alwaysR, rFlags} = {d, dFlags};
          end
        6'b001000: begin // Infinity
            rFlags[ZERO] = 1;
            alwaysR = {d[NEXP+NSIG], {NEXP+NSIG{1'b0}}};
          end
        6'b000100: begin // Zero
            si = ra[roundTowardZero] |
                (ra[roundTowardPositive] & ~d[NEXP+NSIG]) |
                (ra[roundTowardNegative] &  d[NEXP+NSIG]);
            alwaysR = {d[NEXP+NSIG], {NEXP-1{1'b1}}, ~si, {NSIG{si}}};
            rFlags[INFINITY] = ~si;
            rFlags[NORMAL]   =  si;
            exception[DIVIDEBYZERO] = 1;
          end
        default: begin : Normal  // Normal and Subnormal
            reg [1:-(2*NSIG+1)] xa[CLOG2_NSIG:1], xb[CLOG2_NSIG:1];
            reg [2:-(3*NSIG+2)] x[CLOG2_NSIG:0];

            x[0] = 0;
            x[0][0:-(NSIG+1)] = x0;

            for(i = 0; i < CLOG2_NSIG; i = i + 1)
              begin
                // Iteration i
                xa[i+1] = dSigWire * x[i][0:-(NSIG+1)]; // D*xi
                xb[i+1] = (2 << (2*NSIG+1)) - xa[i+1];  // 2 - D*xi
                x[i+1]  = xb[i+1] * x[i][0:-(NSIG+1)];  // (2 - D*xi) * xi
              end
            
            rExp = -dExp;
            
            sigIn = x[CLOG2_NSIG][0:-(3*NSIG+2)] << ~x[CLOG2_NSIG][0];
            normExp[0] = ~x[CLOG2_NSIG][0];
            expIn = rExp - normExp;
            
            if (~|sigOut)
              begin
                rFlags[ZERO] = 1;
                alwaysR = {ra[roundTowardNegative], {NEXP+NSIG{1'b0}}};
              end
            else if (expOut < EMIN)
              begin
                rFlags[SUBNORMAL] = 1;
                alwaysR = {d[NEXP+NSIG], {NEXP{1'b0}}, sigOut[0:1-NSIG]};
              end
            else if (expOut > EMAX)
              begin
                si = ra[roundTowardZero] |
                    (ra[roundTowardPositive] & ~d[NEXP+NSIG]) |
                    (ra[roundTowardNegative] &  d[NEXP+NSIG]);
                alwaysR = {d[NEXP+NSIG], {NEXP-1{1'b1}}, ~si, {NSIG{si}}};
                rFlags[INFINITY] = ~si;
                rFlags[NORMAL]   =  si;
                exception[OVERFLOW] = 1;
              end
            else
              begin
                rFlags[NORMAL] = 1;
                rExp = expOut + BIAS;
                alwaysR = {d[NEXP+NSIG], rExp[NEXP-1:0], sigOut[-1:-NSIG]};
              end

            exception[INEXACT] = inexact;
          end
      endcase
    end

  round #(3*NSIG+3,NEXP,NSIG) U1(d[NEXP+NSIG], expIn, sigIn, ra, expOut, sigOut, inexact);

  assign r = alwaysR;
endmodule
