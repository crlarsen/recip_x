`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Copyright: Chris Larsen, 2022
//
// Create Date: 11/07/2022 09:27:02 AM
// Design Name:
// Module Name: recip_x
// Project Name:
// Target Devices:
// Tool Versions:
// Description: Module to compute the reciprocal of a number D.
//              Normally, we want to compute the reciprocal of a divisor so
//              we can avoid floating point division; multiplication by the
//              reciprocal is almost always much faster. And when performing
//              linear algebra the same divisor is often used multiple times
//              for operations such as normalizing a vector.
//
//              In its present form the module is combinatorial logic.
//              Eventually it will need to be a state machine.
//
//              Inputs:
//              - d: The divisor for which we wish to compute the reciprocal.
//              - ra: The rounding attribute to be used when truncating the
//                    result to fit into the final binary16/-32/-64 result.
//              Outputs:
//              - r: The computed reciprocal value.
//              - rFlags: Flags telling the system which type of value (sNaN,
//                qNaN, Infinity, etc.) is being returned by the module.
//              - exception: Exceptions generated by the module.
//
// Dependencies: fp_class.sv
//               ieee-754-flags.vh
//               padder11.v
//               padder24.v
//               PijGij.v
//               round.v
//               X0.v
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module recip_x(d, ra, r, rFlags, exception);
  parameter NEXP = 5;
  parameter NSIG = 10;
  localparam X0WIDTH = 8;
  `include "ieee-754-flags.vh"
  input [NEXP+NSIG:0] d;
  input [NRAS-1:0] ra;
  output [NEXP+NSIG:0] r;
  output [NTYPES-1:0] rFlags;
  reg [NTYPES-1:0] rFlags;
  output [NEXCEPTIONS-1:0] exception;
  reg [NEXCEPTIONS-1:0] exception;

  localparam hNEXP = 5;
  localparam hNSIG = 10;
  localparam sNEXP = 8;
  localparam sNSIG = 23;
  localparam dNEXP = 11;
  localparam dNSIG = 52;
  localparam qNEXP = 15;
  localparam qNSIG = 112;

  wire inexact, inexactH, inexactX;

  wire signed [NEXP+1:0] dExp, expOut, expOutH, expOutX;
  reg signed [NEXP+1:0] rExp, expIn, normExp = 0;
  wire [0:-NSIG] dSigWire, sigOut, sigOutH, sigOutX;
  wire [NTYPES-1:0] dFlags;
  fp_class #(NEXP,NSIG) dClass(d, dExp, dSigWire, dFlags);

  wire [0:-X0WIDTH] x0;
  X0 U0(dSigWire[-1:-hNSIG], x0);

  reg [NSIG+1+2*X0WIDTH+1:0] sigInH;
  reg [0:-(3*NSIG+2)] sigIn;

  reg [NEXP+NSIG:0] alwaysR;

  reg si;
  always @(*)
    begin
      rFlags = 0;
      exception = 0;

      case (dFlags)
        6'b100000: begin // sNaN
            {alwaysR, rFlags} = {d, dFlags};
          end
        6'b010000: begin // qNaN
            {alwaysR, rFlags} = {d, dFlags};
          end
        6'b001000: begin // Infinity
            rFlags[ZERO] = 1;
            alwaysR = {d[NEXP+NSIG], {NEXP+NSIG{1'b0}}};
          end
        6'b000100: begin // Zero
            si = ra[roundTowardZero] |
                (ra[roundTowardPositive] & ~d[NEXP+NSIG]) |
                (ra[roundTowardNegative] &  d[NEXP+NSIG]);
            alwaysR = {d[NEXP+NSIG], {NEXP-1{1'b1}}, ~si, {NSIG{si}}};
            rFlags[INFINITY] = ~si;
            rFlags[NORMAL]   =  si;
            exception[DIVIDEBYZERO] = 1;
          end
        default: begin : Normal  // Normal and Subnormal
            reg [1:-NSIG-X0WIDTH] x1a, x1b;
            reg [2:-NSIG-2*X0WIDTH] x1;

            // Iteration 1
            x1a = dSigWire * x0;                   // D*x0
            x1b = (2 << (NSIG+X0WIDTH)) - x1a;     // 2 - D*x0
            x1 = x1b * x0;                         // (2 - D*x0) * x0

            rExp = -dExp;

            if (NEXP == hNEXP)
              begin
                // Normalize x1
                sigInH = x1 << ~x1[0];
                normExp[0] = ~x1[0];
                expIn = rExp - normExp;
              end
            else
              begin : BINARY32
                reg [1:-(2*NSIG+1)] x2a, x2b;
                reg [2:-(3*NSIG+2)] x2;

                // Iteration 2
                x2a = dSigWire * x1[0:-(NSIG+1)];
                x2b = (2 << (2*NSIG+1)) - x2a;
                x2 = x2b * x1[0:-(NSIG+1)];

                if (NEXP == sNEXP)
                  begin
                    // Normalize x2
                    sigIn = x2[0:-(3*NSIG+2)] << ~x2[0];
                    normExp[0] = ~x2[0];
                    expIn = rExp - normExp;
                  end
                else
                  begin : BINARY64
                    reg [1:-(2*NSIG+1)] x3a, x3b;
                    reg [2:-(3*NSIG+2)] x3;

                    // Iteration 3
                    x3a = dSigWire * x2[0:-(NSIG+1)];
                    x3b = (2 << (2*NSIG+1)) - x3a;
                    x3 = x3b * x2[0:-(NSIG+1)];

                    // Normalize x3
                    sigIn = x3[0:-(3*NSIG+2)] << ~x3[0];
                    normExp[0] = ~x3[0];
                    expIn = rExp - normExp;
                  end
              end

            if (~|sigOut)
              begin
                rFlags[ZERO] = 1;
                alwaysR = {ra[roundTowardNegative], {NEXP+NSIG{1'b0}}};
              end
            else if (expOut < EMIN)
              begin
                rFlags[SUBNORMAL] = 1;
                alwaysR = {d[NEXP+NSIG], {NEXP{1'b0}}, sigOut[0:1-NSIG]};
              end
            else if (expOut > EMAX)
              begin
                si = ra[roundTowardZero] |
                    (ra[roundTowardPositive] & ~d[NEXP+NSIG]) |
                    (ra[roundTowardNegative] &  d[NEXP+NSIG]);
                alwaysR = {d[NEXP+NSIG], {NEXP-1{1'b1}}, ~si, {NSIG{si}}};
                rFlags[INFINITY] = ~si;
                rFlags[NORMAL]   =  si;
                exception[OVERFLOW] = 1;
              end
            else
              begin
                rFlags[NORMAL] = 1;
                rExp = expOut + BIAS;
                alwaysR = {d[NEXP+NSIG], rExp[NEXP-1:0], sigOut[-1:-NSIG]};
              end

            exception[INEXACT]  = inexact;
          end
      endcase
    end

  if (NSIG == hNSIG)
    round #(NSIG+1+2*X0WIDTH,NEXP,NSIG) U1(d[NEXP+NSIG], expIn, sigInH[NSIG+2*X0WIDTH:0], ra, expOutH, sigOutH, inexactH);
  else
    round #(3*NSIG+3,NEXP,NSIG) U1(d[NEXP+NSIG], expIn, sigIn, ra, expOutX, sigOutX, inexactX);
  assign {expOut, sigOut, inexact} = NSIG == hNSIG ? {expOutH, sigOutH, inexactH} : {expOutX, sigOutX, inexactX};

  assign r = alwaysR;
endmodule
